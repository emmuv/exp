BUCK CONVERTER
VS 1 0 DC 110V
VY 1 2 DC 0V;VOLTAGE SOURCE TO MESURE INPUT CURRENT
VG 7 3 PULSE(0V 20V 0 0.1NS 0.1NS 27.28US 50US)
RB 7 6 250
LE 3 4 681.82UH
CE 4 0 8.33UF IC=60V;INITIAL VOLTAGE
L 4 8 40.91UH
R 8 5 3
VX 5 0 DC 0
DM 0 3 DMOD
.MODEL DMOD D(IS=2.2E-15 BV=1800V TT=0)
Q1 2 6 3 QMOD
.MODEL QMOD NPN(IS=6.734F BF=416.4 BR=0.7371 CJC=3.638P CJE=4.493P TR=239.5N TF=301.2P)
.TRAN 1US 1.6MS 1.5MS 1US UIC
.PROBE
.OPTIONS ABSTOL=1N RELTOL=0.01 VNTOL=0.1 ITL5=50000
.FOUR 20KHZ I(VY)
.END